module FP_Cmp();

endmodule