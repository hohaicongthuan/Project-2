module FP_Mul(in_numA, in_numB, out_result);
    parameter DATA_WIDTH = 64;
    parameter EXP_WIDTH = 11;
    parameter MANT_WIDTH = 52;

    input   [DATA_WIDTH - 1:0] in_numA, in_numB;
    output  [DATA_WIDTH - 1:0] out_result;

    wire    result_sign;
    wire    [EXP_WIDTH - 1:0] result_exp, normalised_exp;
    wire    [MANT_WIDTH - 1:0] normalised_mant;
    wire    [105:0] product_mant;

    assign result_sign = in_numA[63] ^ in_numB[63];
    assign result_exp = (normalised_mant == 0) ? 0 : normalised_exp + 1023;
    assign out_result = {result_sign, result_exp, normalised_mant};

    Mant_Mult Mant_Mult_Inst0(
        .in_multiplicand({54'd1, in_numA[51:0]}),
        .in_multiplier({1'b1, in_numB[51:0]}),
        .out_product(product_mant)
    );
    MultNorm MultNorm_Inst0(
        .in_Exp((in_numA[62:52] - 1023) + (in_numB[62:52] - 1023)),
        .in_Mant(product_mant),
        .out_Exp(normalised_exp),
        .out_Mant(normalised_mant)
    );
endmodule