// This module performs sign injection on a given number
// (Normal sign injection, negated sign injection, and XOR-ed sign injection).

module FP_SGNJ();

endmodule