// Data Memory used for testbench

module DMem();

endmodule