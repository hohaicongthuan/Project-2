module ControlUnit();

endmodule