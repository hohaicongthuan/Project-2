module FP_Div();

endmodule