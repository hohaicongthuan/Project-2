// This module compares two given numbers and returns 1 if the result is true
// otherwise, returns 0

module FP_Cmp(in_numA, in_numB, out_data, in_ctrl);
    parameter DATA_WIDTH = 64;

endmodule