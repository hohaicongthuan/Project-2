module FP_AddSub();

endmodule