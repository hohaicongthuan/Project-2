module FP_Mul();

endmodule