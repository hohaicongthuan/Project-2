// Data Memory used for testbench

module DMem(in_data, in_addr, in_wr_en, out_data);

endmodule