module Testbench();

endmodule