module RV64ID_top();

endmodule