module FP_Convert();

endmodule