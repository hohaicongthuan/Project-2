module FP_MinMax();

endmodule