module RV64IMF();

endmodule