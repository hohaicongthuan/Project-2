module RV64IFD_top();

endmodule