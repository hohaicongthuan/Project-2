// This module converts integer number to floating-point number
module IntToFP(in_data, in_int_width, in_signed_unsigned, in_fp_width, out_data);
    input   in_signed_unsigned;
    input   [1:0] in_int_width, in_fp_width;
    input   [63:0] in_data;

    output  [63:0] out_data;

    
endmodule