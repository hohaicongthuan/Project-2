// Instruction Memory module used for testbench

module IMem();

endmodule