module FP_SGNJ();

endmodule