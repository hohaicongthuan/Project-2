module FP_Unit();

endmodule