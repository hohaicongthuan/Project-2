// This module is the top-level of the Floating-point Unit

module FP_Unit();

endmodule