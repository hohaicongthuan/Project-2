// Multiplier Normaliser
module MultNorm(in_Exp, in_Mant, out_Exp, out_Mant);
    parameter EXP_WIDTH = 11;
    parameter MANT_WIDTH = 52;

    input [EXP_WIDTH - 1:0] in_Exp;
    input [MANT_WIDTH * 2 + 1:0] in_Mant;

    output [EXP_WIDTH - 1:0] out_Exp;
    output [MANT_WIDTH - 1:0] out_Mant;

    assign out_Exp = (in_Mant[MANT_WIDTH * 2 + 1]) ? (in_Exp + 1) : in_Exp;
    assign out_Mant = (in_Mant[MANT_WIDTH * 2 + 1]) ? in_Mant[MANT_WIDTH * 2:53] : in_Mant[MANT_WIDTH * 2 - 1:52];
endmodule